module frogcell(
	input logic clock, reset,
	input logic l, d, u, r,
	output logic ison
);

endmodule 