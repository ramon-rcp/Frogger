module add10_tb();

	logic [8:0] a;
	logic [8:0] b;
	logic [8:0] s;
	logic c;
	
	add10 dut (.a, .b, .s, .c);
	
	initial begin
		a = 9'b000000000; b = 9'b000001010;
		#100; a = 9'b111111000; b = 9'b000000111;
		#100; a = 9'b100000000; b = 9'b100000000;
		#100; a = 9'b100000000; b = 9'b100000000;
		#100; a = 9'b111110000; b = 9'b000010000;
		#100; a = 9'b011110000; b = 9'b000010000;
		#100; a = 9'b101110000; b = 9'b100010000;
		#100;
		
		$stop;
	end 
	
endmodule 